library ieee;
use ieee.std_logic_1164.all;

entity top__proj__ is
  -- Port declarations
  -- port (
    -- p_i_NAME: in|inout|out std_logic|std_logic_vector();
  -- );
end top__proj__;

architecture arch_top__proj__ of top__proj__ is

  -- Submodule instantiation
  -- component submodule_name
    -- generic (
      -- g_PARAM: type := DEFAULT_VALUE
    -- );
    -- port (
      -- p_i_SUB_NAME: in|inout|out type;
    -- );
  -- end component;

begin

  -- i_submodule_name: submodule_name
    -- generic map (
      -- g_PARAM => VALUE
    -- )
    -- port map (
      -- p_i_SUB_NAME => port|signal,
    -- );

end arch_top__proj__;

