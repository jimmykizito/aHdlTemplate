library ieee;
use ieee.std_logic_1164.all;

--! Module description.
entity top___proj__ is
  -- generic (
    -- _PARAM: type := DEFAULT_VALUE;
  -- );
  -- Port declarations
  -- port (
    -- i|io|o_port_name: in|inout|out type;
  -- );
end entity top___proj__;

architecture rtl of top___proj__ is

  -- Submodule instantiation
  -- component submodule_name
    -- generic (
      -- _PARAM: type := DEFAULT_VALUE;
    -- );
    -- port (
      -- i|io|o_port_name: in|inout|out type;
    -- );
  -- end component;

begin

  -- u_submodule_name: submodule_name
    -- generic map (
      -- _PARAM => VALUE,
    -- )
    -- port map (
      -- i|io|o_port_name => port|signal,
    -- );

end architecture rtl;
