library ieee;
use ieee.std_logic_1164.all;

--! Module description.
entity top___proj__ is
  -- generic (
    -- g_PARAM: type := DEFAULT_VALUE;
  -- );
  -- Port declarations
  -- port (
    -- p_i_NAME: in|inout|out std_logic|std_logic_vector();
  -- );
end top___proj__;

architecture arch_top___proj__ of top___proj__ is

  -- Submodule instantiation
  -- component submodule_name
    -- generic (
      -- g_PARAM: type := DEFAULT_VALUE
    -- );
    -- port (
      -- p_i_SUB_NAME: in|inout|out type;
    -- );
  -- end component;

begin

  -- i_submodule_name: submodule_name
    -- generic map (
      -- g_PARAM => VALUE
    -- )
    -- port map (
      -- p_i_SUB_NAME => port|signal,
    -- );

end arch_top___proj__;
